package cnn_pkg;
  import uvm_pkg::*;

  `include "cnn_sequence_item.sv";
  `include "cnn_sequence.sv";
  `include "cnn_sequencer.sv";
  `include "cnn_driver.sv";
  `include "cnn_monitor.sv";
  `include "cnn_agent.sv";
  `include "cnn_scoreboard.sv";
  `include "cnn_env.sv";
  `include "cnn_test.sv";
endpackage
